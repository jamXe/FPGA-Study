//---------------------------------------------------------------------------
//--	文件名		:	A4_Ked1.v
//--	作者		:	ZIRCON
//--	描述		:	KEY控制LED
//--	修订历史	:	2014-1-1
//---------------------------------------------------------------------------
module A4_Key1				//方法1
(
	//输入端口
	KEY0,KEY1,KEY2,KEY3,KEY4,KEY5,KEY6,KEY7,
	//输出端口
	LED0,LED1,LED2,LED3,LED4,LED5,LED6,LED7
);

//---------------------------------------------------------------------------
//--	外部端口声明
//---------------------------------------------------------------------------
input   KEY0,KEY1,KEY2,KEY3,KEY4,KEY5,KEY6,KEY7;	//对应开发板上的KEY
output  LED0,LED1,LED2,LED3,LED4,LED5,LED6,LED7;	//对应开发板上的LED

//---------------------------------------------------------------------------
//--	逻辑功能实现	
//---------------------------------------------------------------------------	
assign LED0 = KEY0;	//触摸按键1控制D1
assign LED1 = KEY1;	//触摸按键2控制D2
assign LED2 = KEY2;	//触摸按键3控制D3
assign LED3 = KEY3;	//触摸按键4控制D4
assign LED4 = KEY4;	//实体按键1控制D5
assign LED5 = KEY5;	//实体按键2控制D6
assign LED6 = KEY6;	//实体按键3控制D7
assign LED7 = KEY7;	//实体按键4控制D8

endmodule					//模块的结束


//module A4_Mini_Key      	//方法2
//(
//  input  [7:0] KEY,		//输入端口声明
//	 output [7:0] LED    	//输出端口声明
//);
//    
//  assign LED = KEY;  	//8个按键控制8个LED
//    
//endmodule              	//模块的结束