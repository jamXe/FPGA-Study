//---------------------------------------------------------------------------
//--	文件名		:	A4_Vote3.v
//--	作者		:	ZIRCON
//--	描述		:	三人表决器（行为描述方式）
//--	修订历史	:	2014-1-1
//---------------------------------------------------------------------------
module A4_Vote3			//模块名A4_Vote3,即模块的开始
(
	//输入端口
	A,B,C,
	//输出端口
	L
);
//---------------------------------------------------------------------------
//--	外部端口声明
//---------------------------------------------------------------------------
input   		A;          //模块的输入端口A
input   		B;          //模块的输入端口B
input   		C;          //模块的输入端口C
output reg 	L;          //模块的输出端口L

//---------------------------------------------------------------------------
//--	逻辑功能实现	
//---------------------------------------------------------------------------
always @ (A,C,B)			//always在组合逻辑中的用法
begin							//always @ (A,B,C)解析：只要A,B,C
	case({A,B,C})			//其中有一个信号有变化便会执行begin中的case语句
		3'b000: L = 1'b0;	//也可以写成always @ (*)，与always @ (A,B,C)功能相同
		3'b001: L = 1'b0;	//{A,B,C}解析：把A,B,C三条线合成一条总线
		3'b010: L = 1'b0;	//举例说明：{1'b1,1'b0}=2'b10
		3'b011: L = 1'b1;	//
		3'b100: L = 1'b0;
		3'b101: L = 1'b1;
		3'b110: L = 1'b1;
		3'b111: L = 1'b1;
		default:L = 1'bx;	//不要省略
	endcase					//case语句的结束
end							//begin语句的结束

endmodule					//module语句的结束
