//---------------------------------------------------------------------------
//--	文件名		:	A4_Ad_Top.v
//--	作者		:	ZIRCON
//--	描述		:	AD的顶层文件,用于将AD获得的电压值显示到数码管上
//--	修订历史	:	2014-1-1
//---------------------------------------------------------------------------
module A4_Ad_Top
(
	//输入端口
	CLK_50M,RST_N,AD_DATA,
	//输出端口
	AD_CS,AD_CLK,SEG_EN,SEG_DATA		
);

//---------------------------------------------------------------------------
//--	外部端口声明
//---------------------------------------------------------------------------
input					CLK_50M;				//时钟端口,开发板用的50M晶振
input					RST_N;				//复位端口,低电平复位
input					AD_DATA;				//AD数据端口
output				AD_CS;				//AD片选端口
output				AD_CLK;				//AD时钟端口
output	[5:0]		SEG_EN;				//数码管使能端口
output	[7:0]		SEG_DATA;			//数码管数据端口

//---------------------------------------------------------------------------
//--	内部端口声明
//---------------------------------------------------------------------------
wire 		[3:0]		vol_int;				//从A/D转换芯片输出的电压值的整数部分；
wire 		[3:0]		vol_dec;				//从A/D转换芯片输出的电压值的小数部分；

//---------------------------------------------------------------------------
//--	逻辑功能实现	
//---------------------------------------------------------------------------
//例化AD模块
Ad_Module			Ad_Init
(
   .CLK_50M			(CLK_50M			),	//时钟端口
   .RST_N			(RST_N			),	//复位端口
	.AD_CS			(AD_CS			),	//AD片选端口
	.AD_CLK			(AD_CLK			),	//AD时钟，最大不超过1.1MHz
	.AD_DATA			(AD_DATA			),	//AD数据端口
	.o_vol_int		(vol_int			),	//从A/D转换芯片输出的电压值的整数部分；
	.o_vol_dec		(vol_dec			)	//从A/D转换芯片输出的电压值的小数部分；
);	

//例化数码管
Segled_Module		Segled_Init
(
	.CLK_50M			(CLK_50M			),	//复位端口
	.RST_N			(RST_N			),	//时钟端口
	.SEG_EN			(SEG_EN			),	//数码管使能端口
	.SEG_DATA		(SEG_DATA		),	//数码管数据端口
	.i_vol_int		(vol_int			),	//从A/D转换芯片输出的电压值的整数部分；
	.i_vol_dec		(vol_dec			)	//从A/D转换芯片输出的电压值的小数部分；
);


endmodule
