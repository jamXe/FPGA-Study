//---------------------------------------------------------------------------
//--	文件名		:	A4_Vote2.v
//--	作者		:	ZIRCON
//--	描述		:	三人表决器（数据流描述方式）
//--	修订历史	:	2014-1-1
//---------------------------------------------------------------------------
module A4_Vote2	//模块名A4_Vote2,即模块的开始
(
	//输出端口
	A,B,C,
	//输入端口
	L
);
//---------------------------------------------------------------------------
//--	外部端口声明
//---------------------------------------------------------------------------
input   A;			//模块的输入端口A
input   B;			//模块的输入端口B
input   C;			//模块的输入端口C
output  L;			//模块的输出端口L

//---------------------------------------------------------------------------
//--	逻辑功能实现	
//---------------------------------------------------------------------------
assign L = (B && C) || (A && C) || (A && B);

endmodule			//模块的结束

