//---------------------------------------------------------------------------
//--	文件名		:	A4_Led1.v
//--	作者		:	ZIRCON
//--	描述		:	点亮LED
//--	修订历史	:	2014-1-1
//---------------------------------------------------------------------------
module A4_Led1				//方法1，模块的开始
(	
	//输出端口
	LED0,LED1,LED2,LED3,LED4,LED5,LED6,LED7
);

//---------------------------------------------------------------------------
//--	外部端口声明
//---------------------------------------------------------------------------
output	LED0,LED1,LED2,LED3,LED4,LED5,LED6,LED7;
	
//---------------------------------------------------------------------------
//--	逻辑功能实现	
//---------------------------------------------------------------------------
assign LED0 = 1'b1;	//给LED0端口赋值1'b0,相信有不少读者会对1'b0感兴趣
assign LED1 = 1'b0;	//为什么要写1'b0,不直接写0，
assign LED2 = 1'b0;	//1'b0是指用的1位二进制，而0则等于32'd0，
assign LED3 = 1'b0;	//只有数字没有进制默认就为十进制，并且位宽默认为32位，
assign LED4 = 1'b1;	//尽管1'b0和32'd0结果是相同的，
assign LED5 = 1'b0;	//但是用十进制表示的话会浪费资源，
assign LED6 = 1'b0;	//因为我们的资源是有限的，
assign LED7 = 1'b0;	//所以节约资源从细节做起，养成良好的编程习惯。
	
endmodule					//模块的结束

//module A4_Led1		//方法2，模块的开始
//(
//	LED					//输出端口的声明
//);
//	output	[7:0] LED;	
//	//LED[0]=1'b1,LED[1]=1'b0,LED[2]=1'b0,LED[3]=1'b0,
//	//LED[4]=1'b1,LED[5]=1'b0,LED[6]=1'b0,LED[7]=1'b0,
//	assign LED = 8'b0001_0001;  
//    
//endmodule				//模块的结束
//
//这里要注意的是，不同的方法，管脚分配名称也是不一样的