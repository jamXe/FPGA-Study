//---------------------------------------------------------------------------
//--	文件名		:	A4_Da_Top.v
//--	作者		:	ZIRCON
//--	描述		:	DA的顶层文件,生成频率1KHz的正弦波
//--	修订历史	:	2014-1-1
//---------------------------------------------------------------------------
module A4_Da_Top
(
	//输入端口
	CLK_50M,RST_N,
	//输出端口
	DA_CLK,DA_CS,DA_DIN
);
 
//---------------------------------------------------------------------------
//--	外部端口声明
//---------------------------------------------------------------------------
input 				CLK_50M;				//时钟端口,开发板用的50M晶振	
input 				RST_N;				//复位端口,低电平复位
output 				DA_CLK;				//DA时钟端口
output 				DA_CS;				//DA片选端口
output 				DA_DIN;				//DA数据输出端口
		
//---------------------------------------------------------------------------
//--	内部端口声明
//---------------------------------------------------------------------------
wire		[9:0]		da_data;				//从ROM中读出的DA数据
wire					da_start;			//DA模块的开始标志位

//---------------------------------------------------------------------------
//--	逻辑功能实现	
//---------------------------------------------------------------------------
//例化DA模块
Da_Module	 		Da_Init
(
	.CLK_50M			(CLK_50M			),	//时钟端口,开发板用的50M晶振	
	.RST_N			(RST_N			),	//复位端口,低电平复位
	.DA_CLK			(DA_CLK			),	//DA时钟端口
	.DA_DIN			(DA_DIN			),	//DA数据输出端口
	.DA_CS			(DA_CS			),	//DA片选端口
	.DA_DATA			(da_data			),	//从ROM中读出的DA数据输入给DA模块
	.send_start		(da_start		)	//DA模块的开始标志位
);

//例化DA数据生成模块
Da_Data_Module		Da_Data_Init
(
	.CLK_50M			(CLK_50M			),	//时钟端口,开发板用的50M晶振	
	.RST_N			(RST_N			),	//复位端口,低电平复位
	.da_data			(da_data			),	//从ROM中读出的DA数据
	.da_start		(da_start		)	//DA模块的开始标志位
);

endmodule
 