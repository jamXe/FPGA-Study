//---------------------------------------------------------------------------
//--	文件名		:	A4_Led3.v
//--	作者		:	ZIRCON
//--	描述		:	同样使LED闪烁和之前不同的代码风格
//--	修订历史	:	2014-1-1
//---------------------------------------------------------------------------
module A4_Led3									
(
	//输入端口
	CLK_50M,RST_N,
	//输出端口
	LED1
);
	
//---------------------------------------------------------------------------
//--	外部端口声明
//---------------------------------------------------------------------------
input 			CLK_50M;						//时钟的端口,开发板用的50M晶振
input				RST_N;						//复位的端口,低电平复位
output 			LED1;							//对应开发板上的LED

//---------------------------------------------------------------------------
//--	内部端口声明
//---------------------------------------------------------------------------
reg			 	led_reg;						//定义显示寄存器
reg	[26:0]	time_cnt;					//定义定时寄存器


//设置定时器的时间为1s,计算方法为  (1*10^9)ns / (1/50)ns  50MHz为开发板晶振
parameter SET_TIME_1S = 27'd50_000_000;

//---------------------------------------------------------------------------
//--	逻辑功能实现	
//---------------------------------------------------------------------------
always @ (posedge CLK_50M or negedge RST_N)
	begin
		if(!RST_N)								//判断复位
			begin 		
				led_reg <= 1'b0;				//初始化led_reg值
			end
		else if (time_cnt == SET_TIME_1S)//判断1s时间
			begin
				led_reg <= ~led_reg;			//如果到达1s,显示寄存器将会被取反
				time_cnt <= 1'b0;				//如果到达1s,定时计数器将会被清零
			end
		else time_cnt <= time_cnt + 1'b1;//如果未到1s,定时计数器将会继续累加
	end

assign LED1 = led_reg;						//最后,将显示寄存器的值赋值给端口LED1

endmodule

