//---------------------------------------------------------------------------
//--	文件名		:	A4_Ir_Top.v
//--	作者		:	ZIRCON
//--	描述		:	通过红外遥控器获得信号值并驱动数码管显示
//--	修订历史	:	2014-1-1
//---------------------------------------------------------------------------
module A4_Ir_Top
(
	//输入端口
	CLK_50M,RST_N,IR_DATA,
	//输出端口
	BEEP		
);

//---------------------------------------------------------------------------
//--	外部端口声明
//---------------------------------------------------------------------------
input					CLK_50M;			//时钟的端口,开发板用的50M晶振
input					RST_N;			//复位的端口,低电平复位
input					IR_DATA;			//红外端口
output				BEEP;				//蜂鸣器端口

//---------------------------------------------------------------------------
//--	内部端口声明
//---------------------------------------------------------------------------
wire 		[7:0]		o_ir_data;		//接收到红外的完整数据

//---------------------------------------------------------------------------
//--	逻辑功能实现	
//---------------------------------------------------------------------------
//例化红外模块
Ir_Module			Ir_Module_Init
(
	.CLK_50M			(CLK_50M		),	//时钟端口
	.RST_N			(RST_N		),	//复位端口
	.IR_DATA			(IR_DATA		),	//红外端口
	.o_ir_data		(o_ir_data	)	//接收的红外的完整数据
);	

//例化蜂鸣器模块
Beep_Module			Beep_Init
(
	.CLK_50M			(CLK_50M		),	//时钟端口
	.RST_N			(RST_N		),	//复位端口
	.BEEP				(BEEP			),	//蜂鸣器端口
	.KEY				(o_ir_data	)	//将接收的数据输出给蜂鸣器模块
);

endmodule


