//---------------------------------------------------------------------------
//--	文件名		:	A4_Vote.v
//--	作者		:	ZIRCON
//--	描述		:	三人表决器（结构化描述方式）
//--	修订历史	:	2014-1-1
//---------------------------------------------------------------------------
module A4_Vote1			//模块名A4_Vote1,即模块的开始,方法1
(
	//输入端口
	A,B,C,
	//输出端口
	L
);

//---------------------------------------------------------------------------
//--	外部端口声明
//---------------------------------------------------------------------------
input   A;              //模块的输入端口A
input   B;              //模块的输入端口B
input   C;              //模块的输入端口C
output  L;              //模块的输出端口L

//---------------------------------------------------------------------------
//--	内部端口声明
//---------------------------------------------------------------------------
wire AB,BC,AC;          //内部信号声明AB,BC,AC
	
//---------------------------------------------------------------------------
//--	逻辑功能实现	
//---------------------------------------------------------------------------
and U1(AB,A,B);         //与门（A,B信号进入）（A与B信号即AB输出）          
and U2(BC,B,C);         //与门 同上
and U3(AC,A,C);         //与门 同上
  
or  U4(L,AB,BC,AC);     //或门 同上
     
endmodule					//模块的结束

//module A4_Vote1(A,B,C,L);//模块名A4_Vote1,即模块的开始,方法2
//
////---端口说明 ---------- 
//
//    input   A;					//模块的输入端口A
//    input   B;					//模块的输入端口B
//    input   C;					//模块的输入端口C
//    output  L;					//模块的输出端口L
//
//   wire NAB,NBC,NAC;			//内部信号声明NAB,NBC,NAC（N代表非、取反）
//      
////---功能描述（门级描述方式）---------- 
//      
//   nand U1(NAB,A,B);			//与非门（A,B信号进入）（A与B信号取非、取反即NAB输出）           
//   nand U2(NBC,B,C);			//与非门 同上
//   nand U3(NAC,A,C);			//与非门 同上
//   
//   nand U4(L,NAB,NBC,NAC);	//与非门 同上
//   
//endmodule							//模块的结束
